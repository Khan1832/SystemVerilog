`include "mem_intf.sv"
`include "apb_common.sv"
`include "memory.v"
`include "mem_assert.v"
`include "apb_tx.sv"
`include "apb_gen.sv"
`include "apb_bfm.sv"
`include "apb_mon.sv"
`include "mem_cov.sv"
`include "apb_agent.sv"
`include "mem_sbd.sv"
`include "apb_env.sv"
`include "top.sv"
